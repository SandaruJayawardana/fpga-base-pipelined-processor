module instuction_mem(data_in,data_out,addr,clk,write_en);
	output [15:0] data_out;
	input [15:0] data_in;
	input [9:0] addr;
	input clk,write_en;
	wire [15:0] data_in,data_out;
	wire clk,write_en;
	wire [9:0] addr;
	reg  [15:0] mem [1023:0];
	
	initial 
		begin // Downsampling instructions are Included 
		mem[ 0 ]= 16'b 0000000000000000 ;
		mem[ 1 ]= 16'b 1111000000000000 ;
		mem[ 2 ]= 16'b 0000000000000000 ;
		mem[ 3 ]= 16'b 1101000000000000 ;
		mem[ 4 ]= 16'b 0000000000000000 ;
		mem[ 5 ]= 16'b 1001100110010000 ;
		mem[ 6 ]= 16'b 0000000001111110 ;
		mem[ 7 ]= 16'b 1001101110110000 ;
		mem[ 8 ]= 16'b 1111111000000000 ;
		mem[ 9 ]= 16'b 1001010101010000 ;
		mem[ 10 ]= 16'b 0000000011111101 ;
		mem[ 11 ]= 16'b 1001011101110000 ;
		mem[ 12 ]= 16'b 0000000000000010 ;
		mem[ 13 ]= 16'b 1001100010000000 ;
		mem[ 14 ]= 16'b 0000000000010000 ;
		mem[ 15 ]= 16'b 1001110011000000 ;
		mem[ 16 ]= 16'b 1111111000000001 ;
		mem[ 17 ]= 16'b 1011000000000000 ;
		mem[ 18 ]= 16'b 0000000000000000 ;
		mem[ 19 ]= 16'b 1110001100010000 ;
		mem[ 20 ]= 16'b 1100000000000000 ;
		mem[ 21 ]= 16'b 1011000000000000 ;
		mem[ 22 ]= 16'b 0000000000000000 ;
		mem[ 23 ]= 16'b 1110010000010000 ;
		mem[ 24 ]= 16'b 1100000000000000 ;
		mem[ 25 ]= 16'b 1011000000000000 ;
		mem[ 26 ]= 16'b 0000000000000000 ;
		mem[ 27 ]= 16'b 0001001100110001 ;
		mem[ 28 ]= 16'b 0001000000000101 ;
		mem[ 29 ]= 16'b 1011000000000000 ;
		mem[ 30 ]= 16'b 0000000000000000 ;
		mem[ 31 ]= 16'b 0001010001000001 ;
		mem[ 32 ]= 16'b 1100000000000000 ;
		mem[ 33 ]= 16'b 1011000000000000 ;
		mem[ 34 ]= 16'b 0000000000000000 ;
		mem[ 35 ]= 16'b 1110011000010000 ;
		mem[ 36 ]= 16'b 1100000000000000 ;
		mem[ 37 ]= 16'b 1011000000000000 ;
		mem[ 38 ]= 16'b 0000000000000000 ;
		mem[ 39 ]= 16'b 0001010001000001 ;
		mem[ 40 ]= 16'b 0001000000000101 ;
		mem[ 41 ]= 16'b 0100011001100111 ;
		mem[ 42 ]= 16'b 1011000000000000 ;
		mem[ 43 ]= 16'b 0100011001100111 ;
		mem[ 44 ]= 16'b 0001001100110001 ;
		mem[ 45 ]= 16'b 1100000000000000 ;
		mem[ 46 ]= 16'b 1011000000000000 ;
		mem[ 47 ]= 16'b 0000000000000000 ;
		mem[ 48 ]= 16'b 0001010001000001 ;
		mem[ 49 ]= 16'b 1100000000000000 ;
		mem[ 50 ]= 16'b 1011000000000000 ;
		mem[ 51 ]= 16'b 0000000000000000 ;
		mem[ 52 ]= 16'b 0001001100110001 ;
		mem[ 53 ]= 16'b 0100010001000111 ;
		mem[ 54 ]= 16'b 0001001100110110 ;
		mem[ 55 ]= 16'b 0000000000000000 ;
		mem[ 56 ]= 16'b 0001001100110100 ;
		mem[ 57 ]= 16'b 1110000011000000 ;
		mem[ 58 ]= 16'b 0101001100111000 ;
		mem[ 59 ]= 16'b 0000000000000000 ;
		mem[ 60 ]= 16'b 1110000100110000 ;
		mem[ 61 ]= 16'b 1010000000000000 ;
		mem[ 62 ]= 16'b 1100001000000000 ;
		mem[ 63 ]= 16'b 0011111010101001 ;
		mem[ 64 ]= 16'b 0110000001001000 ;
		mem[ 65 ]= 16'b 0000000000000000 ;
		mem[ 66 ]= 16'b 1001101010100000 ;
		mem[ 67 ]= 16'b 0000000000000001 ;
		mem[ 68 ]= 16'b 0001110111010111 ;
		mem[ 69 ]= 16'b 0000000000000000 ;
		mem[ 70 ]= 16'b 1110000011010000 ;
		mem[ 71 ]= 16'b 0010111011101110 ;
		mem[ 72 ]= 16'b 0110000000010001 ;
		mem[ 73 ]= 16'b 0000000000000000 ;
		mem[ 74 ]= 16'b 1001110111010000 ;
		mem[ 75 ]= 16'b 0000000100000010 ;
		mem[ 76 ]= 16'b 0010101010101010 ;
		mem[ 77 ]= 16'b 1110000011010000 ;
		mem[ 78 ]= 16'b 0011111010111101 ;
		mem[ 79 ]= 16'b 0111000000010001 ;
		mem[ 80 ]= 16'b 0000000000000000 ;
		mem[ 81 ]= 16'b 0000000000000000 ;
		mem[ 82 ]= 16'b 0000000000000000 ;
		mem[ 83 ]= 16'b 1111111100000000 ;
		end
		
	always @(posedge clk)
		begin
			if(write_en==1'b1)
				mem[addr]=data_in;
		end
	assign 	data_out=mem[addr];
endmodule